`ifndef CORETB_H
`define CORETB_H




package CORETB_PACKAGE;

task dg();
begin
   $display("HELLO WORLD!");
 
end 
endtask 


endpackage


`endif